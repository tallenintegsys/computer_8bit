module computer_8bit
/*#(
// Parameter Declarations
parameter <param_name> = <default_value>,
	parameter [<msb>:<lsb>] <param_name> = <default_value>,
	parameter signed [<msb>:<lsb>] <param_name> = <default_value>
	...
)*/

(
	// Input Ports
	input	CLOCK_50,
	input	[3:0]KEY,

	// Output Ports
	output	[17:0]LEDR,
	output	[8:0]LEDG
);

reg phi;
reg res;
reg so;
reg rdy;
reg nmi;
reg irq;
reg [7:0]dbi;
wire [7:0]dbo;
wire rw;
wire sync;
wire [15:0]ab;
wire [7:0]ram_dbi;
wire [7:0]rom_dbi;

clock_divider c_div(CLOCK_50, phi);

address_decode ad(ab, dbi, ram_dbi, rom_dbi, ram_ce, rom_ce);

single_port_rom rom(ab, phi, rom_ce, rom_dbi);

single_port_ram ram(dbo, ab, phi, rw, ram_dbi);

chip_6502 cpu (
	CLOCK_50,    // FPGA clock
	phi,    // 6502 clock
	res,
	so,
	rdy,
	nmi,
	irq,
	dbi,
	dbo,
	rw,
	sync,
	ab);

// The left-hand side of a continuous assignment must be a structural
// net expression.  That is, it must be a net or a concatentation of
// nets, and any index expressions must be constant.

assign	LEDR[15:0] = ab;
assign	LEDG[7:0] = dbo;
assign	res = !KEY[0];

initial begin
	#0
	so = 1;
	rdy = 1;
	nmi = 1;
	irq = 1;
end

// Module Item(s)

endmodule

